module PraticaIV(SW, HEX0, HEX1, HEX2, HEX3, LEDR);
	input [5:0] SW;
	output [0:6] HEX0;
	output [0:6] HEX1;
	output [0:6] HEX2;
	output [0:6] HEX3;
	output [3:0] LEDR;
	
	
endmodule